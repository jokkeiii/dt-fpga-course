`timescale 1ns / 1ps
module NotGate(input a, output y);
  assign y = !a;
endmodule