`timescale 1ns / 1ps

module AndGate(input a, b, output y);
  assign y=a&b;
endmodule
